//----------------------------------------------------------------------
// Copyright (c) 2025 by Niv Weisman
// nw_recorder - typedef for uvm_recorder
//----------------------------------------------------------------------

`ifndef NW_RECORDER_SVH
`define NW_RECORDER_SVH

typedef uvm_recorder nw_recorder;
typedef uvm_tr_database nw_tr_database;
typedef uvm_text_tr_database nw_text_tr_database;
typedef uvm_tr_stream nw_tr_stream;
typedef uvm_text_tr_stream nw_text_tr_stream;

`endif // NW_RECORDER_SVH

//----------------------------------------------------------------------
// Copyright (c) 2025 by Niv Weisman
// nw_object - typedef for uvm_object
//----------------------------------------------------------------------

`ifndef NW_OBJECT_SVH
`define NW_OBJECT_SVH

typedef uvm_object nw_object;
typedef uvm_void nw_void;
typedef uvm_status_container nw_status_container;
typedef uvm_copy_map nw_copy_map;
typedef uvm_comparer_options nw_comparer_options;
typedef uvm_packer_options nw_packer_options;
typedef uvm_recorder_options nw_recorder_options;
typedef uvm_printer_knobs nw_printer_knobs;
typedef uvm_scope_stack nw_scope_stack;
typedef uvm_objection nw_objection;
typedef uvm_callbacks_objection nw_callbacks_objection;

`endif // NW_OBJECT_SVH

//----------------------------------------------------------------------
// Copyright (c) 2025 by Niv Weisman
// nw_packer - typedef for uvm_packer
//----------------------------------------------------------------------

`ifndef NW_PACKER_SVH
`define NW_PACKER_SVH

typedef uvm_packer nw_packer;

`endif // NW_PACKER_SVH

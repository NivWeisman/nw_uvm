//----------------------------------------------------------------------
// Copyright (c) 2025 by Niv Weisman
// nw_printer - typedef for uvm_printer
//----------------------------------------------------------------------

`ifndef NW_PRINTER_SVH
`define NW_PRINTER_SVH

typedef uvm_printer nw_printer;
typedef uvm_table_printer nw_table_printer;
typedef uvm_tree_printer nw_tree_printer;
typedef uvm_line_printer nw_line_printer;
typedef uvm_hier_printer_knobs nw_hier_printer_knobs;

`endif // NW_PRINTER_SVH

//----------------------------------------------------------------------
// Copyright (c) 2025 by Niv Weisman
// nw_comparer - typedef for uvm_comparer
//----------------------------------------------------------------------

`ifndef NW_COMPARER_SVH
`define NW_COMPARER_SVH

typedef uvm_comparer nw_comparer;

`endif // NW_COMPARER_SVH

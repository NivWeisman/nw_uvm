//----------------------------------------------------------------------
// Copyright (c) 2025 by Niv Weisman
// nw_root - typedef for uvm_root
//----------------------------------------------------------------------

`ifndef NW_ROOT_SVH
`define NW_ROOT_SVH

typedef uvm_root nw_root;
typedef uvm_top nw_top;
typedef uvm_test_done_objection nw_test_done_objection;

`endif // NW_ROOT_SVH
